/*
# KERNEL: UVM_INFO @ 0: reporter [RNTST] Running test my_test...
# KERNEL: UVM_WARNING /home/runner/my_testbench_pkg.svh(79) @ 10: uvm_test_top [] Hello World!
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 10: reporter [FIFO] wdata =   x rdata =   x wfull = 0 rempty = 1 winc = x rinc = x
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 30: reporter [FIFO] wdata =   x rdata =   x wfull = 0 rempty = 1 winc = x rinc = x
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 50: reporter [FIFO] wdata = 121 rdata =   x wfull = 0 rempty = 1 winc = 1 rinc = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 70: reporter [FIFO] wdata = 230 rdata = 121 wfull = 0 rempty = 1 winc = 1 rinc = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 90: reporter [FIFO] wdata = 192 rdata = 121 wfull = 0 rempty = 1 winc = 1 rinc = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 110: reporter [FIFO] wdata =   7 rdata = 121 wfull = 0 rempty = 1 winc = 1 rinc = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 130: reporter [FIFO] wdata = 187 rdata = 121 wfull = 0 rempty = 1 winc = 1 rinc = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 150: reporter [FIFO] wdata = 220 rdata = 121 wfull = 0 rempty = 1 winc = 1 rinc = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 170: reporter [FIFO] wdata = 106 rdata = 121 wfull = 0 rempty = 1 winc = 1 rinc = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 190: reporter [FIFO] wdata = 101 rdata = 121 wfull = 0 rempty = 1 winc = 1 rinc = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 210: reporter [FIFO] wdata = 205 rdata = 121 wfull = 0 rempty = 1 winc = 1 rinc = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 230: reporter [FIFO] wdata = 162 rdata = 121 wfull = 0 rempty = 1 winc = 1 rinc = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 250: reporter [FIFO] wdata = 228 rdata = 121 wfull = 0 rempty = 0 winc = 1 rinc = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 270: reporter [FIFO] wdata = 147 rdata = 121 wfull = 0 rempty = 0 winc = 1 rinc = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 290: reporter [FIFO] wdata = 175 rdata = 121 wfull = 0 rempty = 0 winc = 1 rinc = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 310: reporter [FIFO] wdata =  56 rdata = 121 wfull = 0 rempty = 0 winc = 1 rinc = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 330: reporter [FIFO] wdata =  46 rdata = 121 wfull = 0 rempty = 0 winc = 1 rinc = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 350: reporter [FIFO] wdata = 145 rdata = 121 wfull = 0 rempty = 0 winc = 1 rinc = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 370: reporter [FIFO] wdata =  97 rdata = 121 wfull = 1 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 390: reporter [FIFO] wdata = 158 rdata = 230 wfull = 1 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 410: reporter [FIFO] wdata =  72 rdata = 230 wfull = 1 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 430: reporter [FIFO] wdata =  95 rdata = 230 wfull = 1 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 450: reporter [FIFO] wdata = 227 rdata = 230 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 470: reporter [FIFO] wdata = 212 rdata = 192 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 490: reporter [FIFO] wdata =  50 rdata = 192 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 510: reporter [FIFO] wdata = 253 rdata = 192 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 530: reporter [FIFO] wdata =  53 rdata =   7 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 550: reporter [FIFO] wdata = 218 rdata =   7 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 570: reporter [FIFO] wdata = 236 rdata =   7 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 590: reporter [FIFO] wdata = 107 rdata =   7 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 610: reporter [FIFO] wdata =  87 rdata = 187 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 630: reporter [FIFO] wdata = 176 rdata = 187 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 650: reporter [FIFO] wdata = 118 rdata = 187 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 670: reporter [FIFO] wdata = 169 rdata = 220 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 690: reporter [FIFO] wdata =  73 rdata = 220 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 710: reporter [FIFO] wdata =  86 rdata = 220 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 730: reporter [FIFO] wdata = 208 rdata = 220 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 750: reporter [FIFO] wdata = 183 rdata = 106 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 770: reporter [FIFO] wdata =  11 rdata = 106 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 790: reporter [FIFO] wdata = 204 rdata = 106 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 810: reporter [FIFO] wdata = 250 rdata = 101 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 830: reporter [FIFO] wdata = 149 rdata = 101 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 850: reporter [FIFO] wdata = 157 rdata = 101 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 870: reporter [FIFO] wdata =  18 rdata = 101 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 890: reporter [FIFO] wdata = 244 rdata = 205 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 910: reporter [FIFO] wdata =  67 rdata = 205 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 930: reporter [FIFO] wdata = 255 rdata = 205 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 950: reporter [FIFO] wdata =  40 rdata = 162 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 970: reporter [FIFO] wdata = 190 rdata = 162 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 990: reporter [FIFO] wdata = 193 rdata = 162 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1010: reporter [FIFO] wdata =  49 rdata = 162 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1030: reporter [FIFO] wdata =  14 rdata = 228 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1050: reporter [FIFO] wdata =  88 rdata = 228 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1070: reporter [FIFO] wdata =  15 rdata = 228 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1090: reporter [FIFO] wdata =  51 rdata = 147 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1110: reporter [FIFO] wdata = 196 rdata = 147 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1130: reporter [FIFO] wdata = 194 rdata = 147 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1150: reporter [FIFO] wdata =  45 rdata = 147 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1170: reporter [FIFO] wdata =   5 rdata = 175 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1190: reporter [FIFO] wdata =  74 rdata = 175 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1210: reporter [FIFO] wdata = 252 rdata = 175 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1230: reporter [FIFO] wdata =  27 rdata =  56 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1250: reporter [FIFO] wdata = 167 rdata =  56 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1270: reporter [FIFO] wdata = 160 rdata =  56 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1290: reporter [FIFO] wdata =   6 rdata =  56 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1310: reporter [FIFO] wdata = 217 rdata =  46 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1330: reporter [FIFO] wdata =  25 rdata =  46 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1350: reporter [FIFO] wdata = 198 rdata =  46 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1370: reporter [FIFO] wdata = 224 rdata = 145 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1390: reporter [FIFO] wdata = 103 rdata = 145 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1410: reporter [FIFO] wdata =  91 rdata = 145 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1430: reporter [FIFO] wdata = 188 rdata = 145 wfull = 0 rempty = 0 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1450: reporter [FIFO] wdata = 138 rdata = 121 wfull = 0 rempty = 1 winc = 0 rinc = 1
# KERNEL: UVM_INFO /home/build/vlib1/vlib/uvm-1.2/src/base/uvm_objection.svh(1271) @ 1450: reporter [TEST_DONE] 'run' phase is ready to proceed to the 'extract' phase
# KERNEL: UVM_INFO /home/build/vlib1/vlib/uvm-1.2/src/base/uvm_report_server.svh(869) @ 1450: reporter [UVM/REPORT/SERVER] 
# KERNEL: --- UVM Report Summary ---
# KERNEL: 
# KERNEL: ** Report counts by severity
# KERNEL: UVM_INFO :   76
# KERNEL: UVM_WARNING :    1
# KERNEL: UVM_ERROR :    0
# KERNEL: UVM_FATAL :    0
# KERNEL: ** Report counts by id
# KERNEL: []     1
# KERNEL: [FIFO]    73
# KERNEL: [RNTST]     1
# KERNEL: [TEST_DONE]     1
# KERNEL: [UVM/RELNOTES]     1
# KERNEL: 
# RUNTIME: Info: RUNTIME_0068 uvm_root.svh (521): $finish called.
# KERNEL: Time: 1450 ns,  Iteration: 62,  Instance: /TestBenchTop,  Process: @INITIAL#42_3@.
# KERNEL: stopped at time: 1450 ns
# VSIM: Simulation has finished. There are no more test vectors to simulate.
# VSIM: Simulation has finished.
Done
*/
interface dut_if  #(parameter DSIZE = 8, parameter ASIZE = 4) (); 

  logic [DSIZE-1:0] rdata; 
	logic wfull; 
	logic rempty; 
	logic [DSIZE-1:0] wdata; 
	logic winc, wclk, wrst_n; 
	logic rinc, rclk, rrst_n; 
	
endinterface: dut_if 

`include "uvm_macros.svh"
`include "my_testbench_pkg.svh"

module TestBenchTop (); 


	import uvm_pkg::*;
	import my_testbench_pkg::*;
	
	dut_if _if(); 
	fifo1 dut(
		.rdata(_if.rdata), 
		.wfull(_if.wfull), 
	    .rempty(_if.rempty), 
      	.wdata(_if.wdata), 
		.winc(_if.winc), .wclk(_if.wclk), .wrst_n(_if.wrst_n), 
		.rinc(_if.rinc), .rclk(_if.rclk), .rrst_n(_if.rrst_n) 
	);
	
	//clock generator 
	initial begin 
		_if.wclk = 0; 
		_if.rclk = 0; 
		fork 
			forever #10ns _if.wclk = ~_if.wclk; 
			forever #35ns _if.rclk = ~_if.rclk; 
		join
	end 
	

	initial begin 
		 // Place the interface into the UVM configuration database
		uvm_config_db#(virtual dut_if)::set(null, "*", "dut_vif", _if);
		run_test("my_test"); 
	end 
	
	initial begin 
		$dumpfile("dump.vcd");
      $dumpvars(0, TestBenchTop);
	end 

endmodule: TestBenchTop
  