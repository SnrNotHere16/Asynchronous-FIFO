module DebouncePEDNormal();
endmodule