/*
# KERNEL: ASDB file was created in location /home/runner/dataset.asdb
# KERNEL: UVM_INFO @ 0: reporter [RNTST] Running test my_test...
# KERNEL: UVM_WARNING /home/runner/my_testbench_pkg.svh(79) @ 10: uvm_test_top [] Hello World!
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 10: reporter [FIFO] wdata =   x rdata =   x wfull = 0 rempty = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 30: reporter [FIFO] wdata =   x rdata =   x wfull = 0 rempty = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 50: reporter [FIFO] wdata = 188 rdata =   x wfull = 0 rempty = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 70: reporter [FIFO] wdata = 243 rdata = 188 wfull = 0 rempty = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 90: reporter [FIFO] wdata =  96 rdata = 188 wfull = 0 rempty = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 110: reporter [FIFO] wdata =   3 rdata = 188 wfull = 0 rempty = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 130: reporter [FIFO] wdata = 221 rdata = 188 wfull = 0 rempty = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 150: reporter [FIFO] wdata = 238 rdata = 188 wfull = 0 rempty = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 170: reporter [FIFO] wdata =  53 rdata = 188 wfull = 0 rempty = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 190: reporter [FIFO] wdata = 178 rdata = 188 wfull = 0 rempty = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 210: reporter [FIFO] wdata = 102 rdata = 188 wfull = 0 rempty = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 230: reporter [FIFO] wdata =  81 rdata = 188 wfull = 0 rempty = 1
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 250: reporter [FIFO] wdata = 114 rdata = 188 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 270: reporter [FIFO] wdata = 201 rdata = 188 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 290: reporter [FIFO] wdata =  87 rdata = 188 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 310: reporter [FIFO] wdata =  28 rdata = 188 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 330: reporter [FIFO] wdata =  23 rdata = 188 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 350: reporter [FIFO] wdata =  72 rdata = 188 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 370: reporter [FIFO] wdata = 176 rdata = 188 wfull = 1 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 390: reporter [FIFO] wdata =  79 rdata = 243 wfull = 1 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 410: reporter [FIFO] wdata =  36 rdata = 243 wfull = 1 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 430: reporter [FIFO] wdata =  47 rdata = 243 wfull = 1 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 450: reporter [FIFO] wdata = 113 rdata = 243 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 470: reporter [FIFO] wdata = 234 rdata =  96 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 490: reporter [FIFO] wdata = 153 rdata =  96 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 510: reporter [FIFO] wdata = 126 rdata =  96 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 530: reporter [FIFO] wdata = 154 rdata =   3 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 550: reporter [FIFO] wdata = 237 rdata =   3 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 570: reporter [FIFO] wdata = 118 rdata =   3 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 590: reporter [FIFO] wdata =  53 rdata =   3 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 610: reporter [FIFO] wdata =  43 rdata = 221 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 630: reporter [FIFO] wdata =  88 rdata = 221 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 650: reporter [FIFO] wdata = 187 rdata = 221 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 670: reporter [FIFO] wdata =  84 rdata = 238 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 690: reporter [FIFO] wdata =  36 rdata = 238 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 710: reporter [FIFO] wdata =  43 rdata = 238 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 730: reporter [FIFO] wdata = 104 rdata = 238 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 750: reporter [FIFO] wdata = 219 rdata =  53 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 770: reporter [FIFO] wdata = 133 rdata =  53 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 790: reporter [FIFO] wdata = 102 rdata =  53 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 810: reporter [FIFO] wdata = 125 rdata = 178 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 830: reporter [FIFO] wdata = 202 rdata = 178 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 850: reporter [FIFO] wdata =  78 rdata = 178 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 870: reporter [FIFO] wdata =   9 rdata = 178 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 890: reporter [FIFO] wdata = 250 rdata = 102 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 910: reporter [FIFO] wdata =  33 rdata = 102 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 930: reporter [FIFO] wdata = 127 rdata = 102 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 950: reporter [FIFO] wdata =  20 rdata =  81 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 970: reporter [FIFO] wdata = 223 rdata =  81 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 990: reporter [FIFO] wdata = 224 rdata =  81 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1010: reporter [FIFO] wdata =  24 rdata =  81 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1030: reporter [FIFO] wdata = 135 rdata = 114 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1050: reporter [FIFO] wdata =  44 rdata = 114 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1070: reporter [FIFO] wdata =   7 rdata = 114 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1090: reporter [FIFO] wdata =  25 rdata = 201 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1110: reporter [FIFO] wdata =  98 rdata = 201 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1130: reporter [FIFO] wdata = 225 rdata = 201 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1150: reporter [FIFO] wdata = 150 rdata = 201 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1170: reporter [FIFO] wdata = 130 rdata =  87 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1190: reporter [FIFO] wdata = 165 rdata =  87 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1210: reporter [FIFO] wdata = 254 rdata =  87 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1230: reporter [FIFO] wdata = 141 rdata =  28 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1250: reporter [FIFO] wdata =  83 rdata =  28 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1270: reporter [FIFO] wdata =  80 rdata =  28 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1290: reporter [FIFO] wdata = 131 rdata =  28 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1310: reporter [FIFO] wdata = 236 rdata =  23 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1330: reporter [FIFO] wdata = 140 rdata =  23 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1350: reporter [FIFO] wdata =  99 rdata =  23 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1370: reporter [FIFO] wdata = 112 rdata =  72 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1390: reporter [FIFO] wdata = 179 rdata =  72 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1410: reporter [FIFO] wdata =  45 rdata =  72 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1430: reporter [FIFO] wdata = 222 rdata =  72 wfull = 0 rempty = 0
# KERNEL: UVM_INFO /home/runner/design.sv(223) @ 1450: reporter [FIFO] wdata = 197 rdata = 188 wfull = 0 rempty = 1
# KERNEL: UVM_INFO /home/build/vlib1/vlib/uvm-1.2/src/base/uvm_objection.svh(1271) @ 1450: reporter [TEST_DONE] 'run' phase is ready to proceed to the 'extract' phase
# KERNEL: UVM_INFO /home/build/vlib1/vlib/uvm-1.2/src/base/uvm_report_server.svh(869) @ 1450: reporter [UVM/REPORT/SERVER] 
# KERNEL: --- UVM Report Summary ---
# KERNEL: 
# KERNEL: ** Report counts by severity
# KERNEL: UVM_INFO :   76
# KERNEL: UVM_WARNING :    1
# KERNEL: UVM_ERROR :    0
# KERNEL: UVM_FATAL :    0
# KERNEL: ** Report counts by id
# KERNEL: []     1
# KERNEL: [FIFO]    73
# KERNEL: [RNTST]     1
# KERNEL: [TEST_DONE]     1
# KERNEL: [UVM/RELNOTES]     1
# KERNEL: 
# RUNTIME: Info: RUNTIME_0068 uvm_root.svh (521): $finish called.
# KERNEL: Time: 1450 ns,  Iteration: 62,  Instance: /TestBenchTop,  Process: @INITIAL#42_3@.
# KERNEL: stopped at time: 1450 ns
# VSIM: Simulation has finished. There are no more test vectors to simulate.
# VSIM: Simulation has finished.
Done
*/
interface dut_if  #(parameter DSIZE = 8, parameter ASIZE = 4) (); 

  logic [DSIZE-1:0] rdata; 
	logic wfull; 
	logic rempty; 
	logic [DSIZE-1:0] wdata; 
	logic winc, wclk, wrst_n; 
	logic rinc, rclk, rrst_n; 
	
endinterface: dut_if 

`include "uvm_macros.svh"
`include "my_testbench_pkg.svh"

module TestBenchTop (); 


	import uvm_pkg::*;
	import my_testbench_pkg::*;
	
	dut_if _if(); 
	fifo1 dut(
		.rdata(_if.rdata), 
		.wfull(_if.wfull), 
	    .rempty(_if.rempty), 
      	.wdata(_if.wdata), 
		.winc(_if.winc), .wclk(_if.wclk), .wrst_n(_if.wrst_n), 
		.rinc(_if.rinc), .rclk(_if.rclk), .rrst_n(_if.rrst_n) 
	);
	
	//clock generator 
	initial begin 
		_if.wclk = 0; 
		_if.rclk = 0; 
		fork 
			forever #10ns _if.wclk = ~_if.wclk; 
			forever #35ns _if.rclk = ~_if.rclk; 
		join
	end 
	

	initial begin 
		 // Place the interface into the UVM configuration database
		uvm_config_db#(virtual dut_if)::set(null, "*", "dut_vif", _if);
		run_test("my_test"); 
	end 
	
	initial begin 
		$dumpfile("dump.vcd");
      $dumpvars(0, TestBenchTop);
	end 

endmodule: TestBenchTop
  