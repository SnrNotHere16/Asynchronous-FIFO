
module TestBenchTop (); 




endmodule: TestBenchTop