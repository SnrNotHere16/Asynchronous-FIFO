module AsynchronousFIFO_dut(); 



endmodule: AsynchronousFIFO_dut